library verilog;
use verilog.vl_types.all;
entity Washing_Machine_States_vlg_vec_tst is
end Washing_Machine_States_vlg_vec_tst;
