library verilog;
use verilog.vl_types.all;
entity LED_dot_matrix_vlg_vec_tst is
end LED_dot_matrix_vlg_vec_tst;
