

//点阵玩一下

module LED_dot_matrix(clk, rst, clr, second, state, H, L);

	input clk, rst, clr;
	reg [13:0] posclk_cnt;
	reg clk_9375;
	
	

	input [2:0] state;
	localparam Free = 3'b000;
	localparam Water_supply = 3'b001;
	localparam Rinsing = 3'b011; //3
	localparam Water_draining = 3'b010;
	localparam Dehydrating = 3'b110;
	localparam Warning = 3'b100;
	
	input second;
	reg flip;
	output reg [15:0] H, L;
	
	localparam Row_1 = 16'b0111_1111_1111_1111;
	localparam Row_2 = 16'b1011_1111_1111_1111;
	localparam Row_3 = 16'b1101_1111_1111_1111;
	localparam Row_4 = 16'b1110_1111_1111_1111;
	localparam Row_5 = 16'b1111_0111_1111_1111;
	localparam Row_6 = 16'b1111_1011_1111_1111;
	localparam Row_7 = 16'b1111_1101_1111_1111;
	localparam Row_8 = 16'b1111_1110_1111_1111;
	localparam Row_9 = 16'b1111_1111_0111_1111;
	localparam Row_10 = 16'b1111_1111_1011_1111;
	localparam Row_11 = 16'b1111_1111_1101_1111;
	localparam Row_12 = 16'b1111_1111_1110_1111;
	localparam Row_13 = 16'b1111_1111_1111_0111;
	localparam Row_14 = 16'b1111_1111_1111_1011;
	localparam Row_15 = 16'b1111_1111_1111_1101;
	localparam Row_16 = 16'b1111_1111_1111_1110;
	
	
	always @(posedge clk or negedge rst or negedge clr)	// 分频; 24MHz = '9375' * 2^8 *10
		begin
			if (!rst)
				begin
					posclk_cnt <= 0;
					clk_9375 <= 1;
				end
			else if (!clr)
				begin
					posclk_cnt <= 0;
					clk_9375 <= 1;
				end
			else if (posclk_cnt == 9375)	//9375
				begin
					posclk_cnt <= 0;
					clk_9375 <= 0;
				end
			else
				begin
					posclk_cnt <= posclk_cnt + 1;
					clk_9375 <= 1;
				end
		end
	
	
	always @(negedge second or negedge rst or negedge clr)
		begin
			if (!rst)
				flip <= 0;
			else if (!clr)
				flip <= 0;
			else
				flip <= !flip;
		end
	
	always @(negedge clk_9375 or negedge rst or negedge clr)	//行扫描
		begin
			if (!rst)
				H <= 16'b0111_1111_1111_1111;
			else if (!clr)
				H <= 16'b0111_1111_1111_1111;
			else
				H <= {H[0],H[15:1]};
		end
	
	always @(negedge clk_9375 or negedge rst or negedge clr )
		begin
			if (!rst)
				L <= 16'b1111_1111_1111_1111;
			else if (!clr)
				L <= 16'b1111_1111_1111_1111;
			else
				begin
					case(state)
						Free:
							begin
								if (!flip)
									case(H)
										Row_1:
											L <= 16'b1111_1011_1101_1111; 
										Row_2:
											L <= 16'b1011_1111_1111_1101;
										Row_3:
											L <= 16'b1110_0000_0000_0111;
										Row_4:
											L <= 16'b1110_1111_1111_0111;
										Row_5:
											L <= 16'b1110_1111_1111_0111;
										Row_6:
											L <= 16'b1010_0000_0000_0101;
										Row_7:
											L <= 16'b1110_1111_1111_0111;
										Row_8:
											L <= 16'b1110_1110_0111_0111;
										Row_9:
											L <= 16'b1010_1101_1011_0101;
										Row_10:
											L <= 16'b1110_1010_0101_0111;
										Row_11:
											L <= 16'b1110_1010_0101_0111;
										Row_12:
											L <= 16'b1010_1101_1011_0101;
										Row_13:
											L <= 16'b1110_1110_0111_0111;
										Row_14:
											L <= 16'b1110_1111_1111_0111;
										Row_15:
											L <= 16'b1010_0000_0000_0101;
										Row_16:
											L <= 16'b1111_1111_1111_1111;
									endcase
								else
									case(H)
										Row_1:
											L <= 16'b0111_1011_1101_1110; 
										Row_2:
											L <= 16'b1011_1111_1111_1101;
										Row_3:
											L <= 16'b1110_0000_0000_0111;
										Row_4:
											L <= 16'b1110_1111_1111_0111;
										Row_5:
											L <= 16'b1110_1111_1111_0111;
										Row_6:
											L <= 16'b0010_0000_0000_0100;
										Row_7:
											L <= 16'b1110_1111_1111_0111;
										Row_8:
											L <= 16'b1110_1110_0111_0111;
										Row_9:
											L <= 16'b0010_1101_1011_0100;
										Row_10:
											L <= 16'b1110_1010_0101_0111;
										Row_11:
											L <= 16'b1110_1010_0101_0111;
										Row_12:
											L <= 16'b0010_1101_1011_0100;
										Row_13:
											L <= 16'b1110_1110_0111_0111;
										Row_14:
											L <= 16'b1110_1111_1111_0111;
										Row_15:
											L <= 16'b1010_0000_0000_0101;
										Row_16:
											L <= 16'b0111_1111_1111_1110;
									endcase
							end
						Water_supply:
							begin
								if (!flip)
									case(H)
										Row_1:
											L <= 16'b1111_1111_1111_1111; 
										Row_2:
											L <= 16'b1111_1100_0011_1111;
										Row_3:
											L <= 16'b1111_0011_1100_1111;
										Row_4:
											L <= 16'b1110_1111_1111_0111;
										Row_5:
											L <= 16'b1101_1111_1111_1011;
										Row_6:
											L <= 16'b1101_1111_1111_1011;
										Row_7:
											L <= 16'b1011_1111_1111_1101;
										Row_8:
											L <= 16'b1011_1111_1111_1101;
										Row_9:
											L <= 16'b1011_1111_1111_1101;
										Row_10:
											L <= 16'b1011_1111_1111_1101;
										Row_11:
											L <= 16'b1101_0011_1100_1011;
										Row_12:
											L <= 16'b1100_1101_1011_0011;
										Row_13:
											L <= 16'b1110_1110_0111_0111;
										Row_14:
											L <= 16'b1111_0011_1100_1111;
										Row_15:
											L <= 16'b1111_1100_0011_1111;
										Row_16:
											L <= 16'b1111_1111_1111_1111;
									endcase
								else
									case(H)
										Row_1:
											L <= 16'b1111_1111_1111_1111; 
										Row_2:
											L <= 16'b1111_1100_0011_1111;
										Row_3:
											L <= 16'b1111_0011_1100_1111;
										Row_4:
											L <= 16'b1110_1111_1111_0111;
										Row_5:
											L <= 16'b1101_0011_1100_1011;
										Row_6:
											L <= 16'b1100_1101_1011_0011;
										Row_7:
											L <= 16'b1011_1110_0111_1101;
										Row_8:
											L <= 16'b1011_1111_1111_1101;
										Row_9:
											L <= 16'b1011_1111_1111_1101;
										Row_10:
											L <= 16'b1011_1111_1111_1101;
										Row_11:
											L <= 16'b1101_1111_1111_1011;
										Row_12:
											L <= 16'b1101_1111_1111_1011;
										Row_13:
											L <= 16'b1110_1111_1111_0111;
										Row_14:
											L <= 16'b1111_0011_1100_1111;
										Row_15:
											L <= 16'b1111_1100_0011_1111;
										Row_16:
											L <= 16'b1111_1111_1111_1111;
									endcase
							end
						Rinsing:
							begin
								if (!flip)
									case(H)
										Row_1:
											L <= 16'b1111_1111_1111_1111; 
										Row_2:
											L <= 16'b1111_1100_0011_1111;
										Row_3:
											L <= 16'b1111_0011_1100_1111;
										Row_4:
											L <= 16'b1110_1111_1111_0111;
										Row_5:
											L <= 16'b1101_1001_1001_1011;
										Row_6:
											L <= 16'b1101_0110_0110_1011;
										Row_7:
											L <= 16'b1011_0111_1110_1101;
										Row_8:
											L <= 16'b1011_0011_1100_1101;
										Row_9:
											L <= 16'b1011_1011_1101_1101;
										Row_10:
											L <= 16'b1011_1011_1101_1101;
										Row_11:
											L <= 16'b1101_1011_1101_1011;
										Row_12:
											L <= 16'b1101_1000_0001_1011;
										Row_13:
											L <= 16'b1110_1111_1111_0111;
										Row_14:
											L <= 16'b1111_0011_1100_1111;
										Row_15:
											L <= 16'b1111_1100_0011_1111;
										Row_16:
											L <= 16'b1111_1111_1111_1111;
									endcase
								else
									case(H)
										Row_1:
											L <= 16'b1111_1111_1111_1111; 
										Row_2:
											L <= 16'b1111_1100_0011_1111;
										Row_3:
											L <= 16'b1111_0011_1100_1111;
										Row_4:
											L <= 16'b1110_1111_1111_0111;
										Row_5:
											L <= 16'b1101_1000_0001_1011;
										Row_6:
											L <= 16'b1101_1101_1011_1011;
										Row_7:
											L <= 16'b1011_1011_1101_1101;
										Row_8:
											L <= 16'b1011_1010_0101_1101;
										Row_9:
											L <= 16'b1011_1010_0101_1101;
										Row_10:
											L <= 16'b1011_1001_1001_1101;
										Row_11:
											L <= 16'b1101_1001_1001_1011;
										Row_12:
											L <= 16'b1101_1001_1001_1011;
										Row_13:
											L <= 16'b1110_1111_1111_0111;
										Row_14:
											L <= 16'b1111_0011_1100_1111;
										Row_15:
											L <= 16'b1111_1100_0011_1111;
										Row_16:
											L <= 16'b1111_1111_1111_1111;
									endcase
							end
						Water_draining:
							begin
								if (!flip)
									case(H)
										Row_1:
											L <= 16'b1111_1111_1111_1111; 
										Row_2:
											L <= 16'b1111_1100_0011_1111;
										Row_3:
											L <= 16'b1111_1110_0111_1111;
										Row_4:
											L <= 16'b1110_0000_0011_1111;
										Row_5:
											L <= 16'b1111_1111_1101_1111;
										Row_6:
											L <= 16'b1110_0001_1101_1111;
										Row_7:
											L <= 16'b1111_1110_1101_1111;
										Row_8:
											L <= 16'b1111_1110_0011_1111;
										Row_9:
											L <= 16'b1111_1111_1111_1111;
										Row_10:
											L <= 16'b1111_1111_0111_1111;
										Row_11:
											L <= 16'b1111_1111_0111_1111;
										Row_12:
											L <= 16'b1111_1110_0011_1111;
										Row_13:
											L <= 16'b1111_1111_1111_1111;
										Row_14:
											L <= 16'b1111_1111_1111_1111;
										Row_15:
											L <= 16'b1111_1111_1111_1111;
										Row_16:
											L <= 16'b1111_1111_1111_1111;
									endcase
								else
									case(H)
										Row_1:
											L <= 16'b1111_1111_1111_1111; 
										Row_2:
											L <= 16'b1111_1100_0011_1111;
										Row_3:
											L <= 16'b1111_1110_0111_1111;
										Row_4:
											L <= 16'b1110_0000_0011_1111;
										Row_5:
											L <= 16'b1111_1111_1101_1111;
										Row_6:
											L <= 16'b1110_0001_1101_1111;
										Row_7:
											L <= 16'b1111_1110_1101_1111;
										Row_8:
											L <= 16'b1111_1110_0011_1111;
										Row_9:
											L <= 16'b1111_1111_1111_1111;
										Row_10:
											L <= 16'b1111_1111_1111_1111;
										Row_11:
											L <= 16'b1111_1111_1111_1111;
										Row_12:
											L <= 16'b1111_1111_1111_1111;
										Row_13:
											L <= 16'b1111_1111_0111_1111;
										Row_14:
											L <= 16'b1111_1111_0111_1111;
										Row_15:
											L <= 16'b1111_1110_0011_1111;
										Row_16:
											L <= 16'b1111_1111_1111_1111;
									endcase
							end
						Dehydrating:
							begin
								if (!flip)
									case(H)
										Row_1:
											L <= 16'b1111_1111_1111_1111; 
										Row_2:
											L <= 16'b1011_1101_1101_1011;
										Row_3:
											L <= 16'b0000_0000_0000_0000;
										Row_4:
											L <= 16'b1011_1101_1101_1011;
										Row_5:
											L <= 16'b1011_1101_1101_1011;
										Row_6:
											L <= 16'b1001_1001_1000_0001;
										Row_7:
											L <= 16'b0110_0110_1101_1011;
										Row_8:
											L <= 16'b0111_1110_1011_1101;
										Row_9:
											L <= 16'b0011_1100_1010_0101;
										Row_10:
											L <= 16'b1011_1101_1010_0101;
										Row_11:
											L <= 16'b1011_1101_1001_1001;
										Row_12:
											L <= 16'b1011_1101_1001_1001;
										Row_13:
											L <= 16'b1000_0001_1001_1001;
										Row_14:
											L <= 16'b1111_1111_1111_1111;
										Row_15:
											L <= 16'b1101_1011_1101_1011;
										Row_16:
											L <= 16'b1101_1011_1101_1011;
									endcase
								else
									case(H)
										Row_1:
											L <= 16'b1111_1111_1111_1111; 
										Row_2:
											L <= 16'b1011_1101_1101_1011;
										Row_3:
											L <= 16'b0000_0000_0000_0000;
										Row_4:
											L <= 16'b1011_1101_1101_1011;
										Row_5:
											L <= 16'b1011_1101_1101_1011;
										Row_6:
											L <= 16'b1001_1001_1000_0001;
										Row_7:
											L <= 16'b0110_0110_1101_1011;
										Row_8:
											L <= 16'b0111_1110_1011_1101;
										Row_9:
											L <= 16'b0011_1100_1010_0101;
										Row_10:
											L <= 16'b1011_1101_1010_0101;
										Row_11:
											L <= 16'b1011_1101_1001_1001;
										Row_12:
											L <= 16'b1011_1101_1001_1001;
										Row_13:
											L <= 16'b1000_0001_1001_1001;
										Row_14:
											L <= 16'b1111_1111_1111_1111;
										Row_15:
											L <= 16'b1011_1101_1011_1101;
										Row_16:
											L <= 16'b1011_1101_1011_1101;
									endcase
							end
						Warning:
							begin
								if (!flip)
									case(H)
										Row_1:
											L <= 16'b1111_1111_1111_1111; 
										Row_2:
											L <= 16'b1111_1110_0111_1111;
										Row_3:
											L <= 16'b1111_1110_0111_1111;
										Row_4:
											L <= 16'b1111_1110_0111_1111;
										Row_5:
											L <= 16'b1101_1110_0111_1011;
										Row_6:
											L <= 16'b1100_1110_0111_0011;
										Row_7:
											L <= 16'b1110_1110_0111_0111;
										Row_8:
											L <= 16'b1111_1110_0111_1111;
										Row_9:
											L <= 16'b1111_1101_1011_1111;
										Row_10:
											L <= 16'b1111_1101_1011_1111;
										Row_11:
											L <= 16'b1111_1101_1011_1111;
										Row_12:
											L <= 16'b1111_1101_1011_1111;
										Row_13:
											L <= 16'b1111_1000_0001_1111;
										Row_14:
											L <= 16'b1100_1110_0111_0011;
										Row_15:
											L <= 16'b1001_1111_1111_1001;
										Row_16:
											L <= 16'b1111_1111_1111_1111;
									endcase
								else
									case(H)
										Row_1:
											L <= 16'b1111_1111_1111_1111; 
										Row_2:
											L <= 16'b1111_1110_0111_1111;
										Row_3:
											L <= 16'b1111_1110_0111_1111;
										Row_4:
											L <= 16'b1111_1110_0111_1111;
										Row_5:
											L <= 16'b1111_1110_0111_1111;
										Row_6:
											L <= 16'b1111_1110_0111_1111;
										Row_7:
											L <= 16'b1111_1110_0111_1111;
										Row_8:
											L <= 16'b1111_1110_0111_1111;
										Row_9:
											L <= 16'b1111_1101_1011_1111;
										Row_10:
											L <= 16'b1001_1101_1011_1001;
										Row_11:
											L <= 16'b1100_1101_1011_0011;
										Row_12:
											L <= 16'b1111_1101_1011_1111;
										Row_13:
											L <= 16'b1111_1000_0001_1111;
										Row_14:
											L <= 16'b1111_1110_0111_1111;
										Row_15:
											L <= 16'b1111_1111_1111_1111;
										Row_16:
											L <= 16'b1111_1111_1111_1111;
									endcase
							end
					endcase
				end
		end
	
endmodule
