library verilog;
use verilog.vl_types.all;
entity Timer_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        clr             : in     vl_logic;
        pause           : in     vl_logic;
        rst             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Timer_vlg_sample_tst;
