library verilog;
use verilog.vl_types.all;
entity Breathing_LED_vlg_vec_tst is
end Breathing_LED_vlg_vec_tst;
